/**
 * \file aes.sv
 * \author Eric Mueller
 * Addapted from aes_starter.sv by bchasnov@hmc.edu, David_Harris@hmc.edu
 */


/* Test AES with cases from FIPS-197 appendix */
module testbench();
   logic clk, load, done, sck, sdi, sdo;
   logic [127:0] key, plaintext, cyphertext, expected;
   logic [255:0] comb;
   logic [8:0]   i;
    
   // device under test
   aes dut(clk, sck, sdi, sdo, load, done);
    
   // test case
   initial begin   
      // Test case from FIPS-197 Appendix A.1, B
      key       <= 128'h2B7E151628AED2A6ABF7158809CF4F3C;
      plaintext <= 128'h3243F6A8885A308D313198A2E0370734;
      expected  <= 128'h3925841D02DC09FBDC118597196A0B32;
      
// Alternate test case from Appendix C.1
//      key       <= 128'h000102030405060708090A0B0C0D0E0F;
//      plaintext <= 128'h00112233445566778899AABBCCDDEEFF;
//      expected  <= 128'h69C4E0D86A7B0430D8CDB78070B4C55A;
   end
    
   // generate clock and load signals
   initial 
     forever begin
        clk = 1'b0; #5;
        clk = 1'b1; #5;
     end
   
   initial begin
      i = 0;
      load = 1'b1;
   end 
   
   assign comb = {plaintext, key};
   // shift in test vectors, wait until done, and shift out result
   always @(posedge clk) begin
      if (i == 256) load = 1'b0;
      if (i<256) begin
         #1; sdi = comb[255-i];
         #1; sck = 1; #5; sck = 0;
         i = i + 1;
      end else if (done && i < 384) begin
         #1; sck = 1; 
         #1; cyphertext[383-i] = sdo;
         #4; sck = 0;
         i = i + 1;
      end else if (i == 384) begin
         if (cyphertext == expected)
           $display("Testbench ran successfully");
         else $display("Error: cyphertext = %h, expected %h",
                       cyphertext, expected);
         $stop();
         
      end
   end   
endmodule


/** 
 * Top level module with SPI interface and SPI core
 * 
 * \param clk    40MHz board clock
 * \param sck    serial clock
 * \param sdi    slave data in, aka MOSI
 * \param sdo    slave data out, aka MISO
 * \param load   load signal from Pi's GPIO pin
 * \param done   done signal to Pi's GPIO pin
 */
module aes(input  logic clk,
           input  logic sck, 
           input  logic sdi,
           output logic sdo,
           input  logic load,
           output logic done);
                    
   logic [127:0]        key, plaintext, cyphertext;
   
   aes_spi spi(sck, sdi, sdo, done, key, plaintext, cyphertext);   
   aes_core core(clk, load, key, plaintext, done, cyphertext);
endmodule


/**
 * SPI interface.  Shifts in key and plaintext Captures ciphertext when done,
 * then shifts it out.
 * 
 * \param sck    serial clock
 * \param sdi    slave data in, aka MOSI
 * \param sdo    slave data out, aka MISO
 * \param done   done signal to Pi's GPIO pin
 * \param key    key read from Pi
 * \param plaintext     plaintext read from Pi
 * \param cyphertext    cyphertext to write back to the Pi
 */
module aes_spi(input  logic sck, 
               input  logic sdi,
               output logic sdo,
               input  logic done,
               output logic [127:0] key, plaintext,
               input  logic [127:0] cyphertext);

   logic                            sdodelayed, wasdone;
   logic [127:0]                    cyphertextcaptured;


   /* Tricky cases to properly change sdo on negedge clk. */

   // assert load
   // apply 256 sclks to shift in key and plaintext, starting with plaintext[0]
   // then deassert load, wait until done
   // then apply 128 sclks to shift out cyphertext, starting with cyphertext[0]
   always_ff @(posedge sck)
     if (!wasdone)  {cyphertextcaptured, plaintext, key} = {cyphertext, plaintext[126:0], key, sdi};
     else           {cyphertextcaptured, plaintext, key} = {cyphertextcaptured[126:0], plaintext, key, sdi}; 
   
   // sdo should change on the negative edge of sck
   always_ff @(negedge sck) begin
      wasdone = done;
      sdodelayed = cyphertextcaptured[126];
   end
    
   // when done is first asserted, shift out msb before clock edge
   assign sdo = (done & !wasdone) ? cyphertext[127] : sdodelayed;
endmodule


/**
 * top level AES encryption module
 * 
 * \param clk          40MHz board clock
 * \param load         raised when encryption should start
 * \param key          key to encrypt
 * \param plaintext    data to encrypt
 * \param done         raised with the encryption is finished
 * \param cyphertext   result of the encryption
 * 
 *   when load is asserted, takes the current key and plaintext
 *   generates cyphertext and asserts done when complete 11 cycles later
 * 
 *   See FIPS-197 with Nk = 4, Nb = 4, Nr = 10
 *
 *   The key and message are 128-bit values packed into an array of 16 bytes as
 *   shown below
 *        [127:120] [95:88] [63:56] [31:24]     S0,0    S0,1    S0,2    S0,3
 *        [119:112] [87:80] [55:48] [23:16]     S1,0    S1,1    S1,2    S1,3
 *        [111:104] [79:72] [47:40] [15:8]      S2,0    S2,1    S2,2    S2,3
 *        [103:96]  [71:64] [39:32] [7:0]       S3,0    S3,1    S3,2    S3,3
 *
 *   Equivalently, the values are packed into four words as given
 *        [127:96]  [95:64] [63:32] [31:0]      w[0]    w[1]    w[2]    w[3]
 */
module aes_core(input  logic         clk, 
                input  logic         load,
                input  logic [127:0] key, 
                input  logic [127:0] plaintext, 
                output logic         done, 
                output logic [127:0] cyphertext);

   /* XXX: write this mofo */
    
endmodule


/**
 * Infamous AES byte substitutions with magic numbers
 * Section 5.1.1, Figure 7
 */
module sbox(input  logic [7:0] a,
            output logic [7:0] y);
            
  // sbox implemented as a ROM
  logic [7:0] sbox[0:255];

  initial   $readmemh("sbox.txt", sbox);
  assign y = sbox[a];
endmodule


/**
 * Even funkier action on columns
 * Section 5.1.3, Figure 9
 * Same operation performed on each of four columns
 */
module mixcolumns(input  logic [127:0] a,
                  output logic [127:0] y);

  mixcolumn mc0(a[127:96], y[127:96]);
  mixcolumn mc1(a[95:64],  y[95:64]);
  mixcolumn mc2(a[63:32],  y[63:32]);
  mixcolumn mc3(a[31:0],   y[31:0]);
endmodule


/**
 * Perform Galois field operations on bytes in a column
 * See EQ(4) from E. Ahmed et al, Lightweight Mix Columns Implementation for AES, AIC09
 * for this hardware implementation
 */
module mixcolumn(input  logic [31:0] a,
                 output logic [31:0] y);
                      
   logic [7:0]       a0, a1, a2, a3, y0, y1, y2, y3, t0, t1, t2, t3, tmp;
        
   assign {a0, a1, a2, a3} = a;
   assign tmp = a0 ^ a1 ^ a2 ^ a3;
    
   galoismult gm0(a0^a1, t0);
   galoismult gm1(a1^a2, t1);
   galoismult gm2(a2^a3, t2);
   galoismult gm3(a3^a0, t3);

   assign y0 = a0 ^ tmp ^ t0;
   assign y1 = a1 ^ tmp ^ t1;
   assign y2 = a2 ^ tmp ^ t2;
   assign y3 = a3 ^ tmp ^ t3;
   assign y = {y0, y1, y2, y3};    
endmodule


/**
 * Multiply by x in GF(2^8) is a left shift
 * followed by an XOR if the result overflows
 * Uses irreducible polynomial x^8+x^4+x^3+x+1 = 00011011
 */
module galoismult(input  logic [7:0] a,
                  output logic [7:0] y);

   logic [7:0]                       ashift;
    
   assign ashift = {a[6:0], 1'b0};
   assign y = a[7] ? (ashift ^ 8'b00011011) : ashift;
endmodule
